Hur man spelar Freeciv

  Ursprungligen av Michael Hohensee (aka Zarchon)

För upplysningar om hur man installerar Freeciv, se INSTALL.sv
För upplysningar om hur man kör Freeciv, se README.sv

Om man aldrig har spelat något av spelen i Civilization-serien
är det bäst om man börjar med att läsa Freecivs handbok som är
tillgänglig vid:

     https://www.freeciv.org/wiki/Manual

För upplysningar om hur man spelar Freeciv, fortsätt läsa!

	När man har fått i gång Freeciv vill man antagligen spela sina
första spel. Man råds att spela ensam några gånger för att få en
känsla för hur saker fungerar, men det är inte nödvändigt. Man kan
lära sig genom att spela mot andra människor eller mot datorn.

Fråga: Vilken är den grundläggande strategin?

	För det första är detta inte en *perfekt* strategi; det är
inte ens en mycket bra strategi. Men låt oss först sätta i gång med att
spela Freeciv. En del av lockelsen hos Freeciv är att utveckla nya
strategier.

	Strategin är indelat i flera steg:

		Det inledande utvidgningsskedet
		Teknologiskt underskede
		Det andra utvidgningsskedet
		Uppbyggnadsskedet
		Den slutgiltiga förintelsen av dina fiender-skedet

Det inledande utvidgningsskedet:

	Detta skede är viktigast. Det första man bör göra är att
grunda städer och utforska sin ö. Man bör ha många städer, mist 7
eller 8.

	Spelets mål är att behärska så många landrutor som möjligt.
När man grundar en stad bör man se till att att dess område inte
kommer att överlappa för mycket med andra städers områden. Man kan se
vilka rutor som används av en stad genom att klicka på den. Kartan
över staden och dess omgivning visar stadens område. Ta hänsyn till
detta och försök samtidigt att hålla dina städer nära varandra. Ju
längre från varandra de är, desto svårare är det att försvara och
förvalta dem i detta skede. (Hänvisning: Försök att grunda städer på
hästar eller nära fisk.)

	När man har 1 eller 2 städer bör man sätta forskningssatsen så
högt som regeringsformen tillåter. Man ska strunta i skattesatsen
eftersom man inte kommer att färdigställa några stadsförbättringar som
kostar underhåll regelbundet. Man bygger i stället bosättare. Varje
stad bör bygga bosättare. Ju fler bosättare man färdigställer, desto
fler städer kan man grunda; ju fler städer man har, desto fortare kan
man forska; ju fortare man kan forska, desto fortare kan man vinna.
När man har fyllt det tillgängliga utrymmet med städer befaller man
sina bosättare att bygga bevattningsanläggningar och vägar.

(Anmärkning: Om matöverskottet i en stad sjunker till +1 på grund
av understöd av för många bosättare och man inte kan flytta om
arbetare så att överskottet blir större låter man staden bygga ett
tempel i stället för bosättare. Om man inte har känner sig hotad av
någon annan spelare än kan man strunta i att bygga krigsenheter ett
tag till.)

	Under denna tid lär man sig teknologier så fort som möjligt.
Det man bör sikta på först är "republik", sedan "folkstyre", sedan
"järnväg", sedan "industrialisering". (Vissa siktar på "monarki" före
"republik".) Så snart som man forskat fram en regeringsform som man
vill använda sätter man i gång en revolution och byter till den nya
regeringsformen när revolutionen är över. Sedan ser man till att
satserna är som man vill ha dem, ty den högsta tillåtna satsen skiljer
sig mellan olika regeringsformer (forskningssatsen sätts så högt som
möjligt av sig själv).

	När man har fått kunskap om folkstyre är man rustad att gå in
i det andra utvidgningsskedet. Det gör man genom att ändra
regeringsform till folkstyre, befalla alla städer att bygga tempel och
sätta överflödssatsen till 100%. När man gör detta börjar alla städer
genast att fira och växer 1 steg varje omgång så länge det finns
matöverskott. När de har blivit tillräckligt stora sätt
överflödssatsen till rimliga 20-40%. Detta försätter dig i det andra
utvidgningsskedet.

	Nackdelen med att sätta överflödssatsen till 100% är att
forskningen avstannar fullständigt. Efter att städerna har vuxit och
forskningssatsen har höjts till ungefär 50% får man åter nya
teknologier, men något saktare. Om man har utforskat ganska mycket
utan att ha hittat någon hotfull motspelare kan det vara bra att
forska så mycket som möjligt tills teknologierna tar för lång tid att
forska fram.

Det andra utvidgningsskedet:

	När städerna har fått en lämplig storlek avvänjer man dem med
överflöd och ökar skattesatsen. När de är nere på ungefär 30% överflöd
ökar man forskningssatsen så mycket man kan utan att skatteinkomsten
blir lägre än utgifterna. När man får järnväg bygger man om alla vägar
till järnvägar, åtminstone alla som är på rutor som används av någon
stads arbetare eller ingår i fjärrvägnätet. (Hänvisning: Utrusta varje
ruta som används av en stad med väg/järnväg. Då gör staden mer nytta.
Det finns ingen anledning att uppgradera mittrutan, den med staden på.
Det görs av sig själv.)

	Nu är det dags att utveckla industrialisering och
krigsteknologier. Man bör börja grunda städer på andra öar och
utforska ordentligt om man inte redan har gjort det. Man bör ta reda
på var fienderna är. Sikta på teknologier som är bra för båtar och
försök färdigställa Magellans Världsomsegling. När man känner dig
beredd går man in i:

Uppbyggnadsskedet:

	Nu bygger man fabriker och kraftverk i städerna. Man försöker
få så hög tillverkningsförmåga som möjligt. Förorening blir ett
problem. Så snart man kan försöker man forska fram masstillverkning
för kollektivtrafik och återvinning för återvinningsanläggning. När
man har gjort alla sina städer till goda tillverkningsanläggningar
bygger man krigsenheter. (Anmärkning: Om man får förbindelse med någon
annan spelare ska man genast bygga några angreppsenheter och minst 1
försvarsenhet för varje stad.)

	När man vill börja angripa någon sätter man forskningssatsen
till 0% och höjer skattesatsen så mycket man kan utan att få upplopp.
Kom ihåg att enheter kan köpas för guld!

Den slutgiltiga förintelsen av dina fiender-skedet:

	Detta kan ske när som helst men det är skojigare med de
framskridna vapnen.

	Välj en förhållandevis svag fiende och skicka över några
båtlaster trupper. Ta över fiendens städer och låt dem bygga fler
enheter för att utplåna resten av fienden. Visa ingen medkänsla!
Intill döden!

Upprepa så ofta som det behövs! ;-)

[Anmärkning för fredliga: Freeciv låter även en spelare vinna genom
att färdigställa och sända iväg ett rymdskepp som anländer till Alfa
Kentauri före alla andra spelares eventuella rymdskepp.]


Ytterligare frågor:

Fråga: Vilka andra strategier finns det?

	Det finns ett antal handledningar och strategianvisningar
tillgängliga vid Freecivs webplats vid:

	 https://www.freeciv.org/wiki/Tutorials

Dessutom beskriver Freecivs inbyggda hjälp en annan strategi.


Fråga: Vilken tidsgräns skall man sätta i flerspelarspel?

	Det beror på antalet spelare. Om man bara är 2 som spelar
klarar man sig vanligtvis med tidsgränsen 0. Om man är > 2 eller en av
de 2 kommer att vara borta från spelet under slumpmässliga tillfällen
och den andre inte vill vänta kan en tidsgräns på 1 minut (när man
sätter tidsgränsen anger man dock tiden i sekunder) vara tillräckligt.
Senare i spelet när det är mer att göra vill man antagligen öka
tidsgränsen till 4 minuter. I allmänhet behövs det längre tid ju fler
spelare man är. Sätt den tidsgräns som passar men kom i håg att det brukar
störa folk om man går över 5 minuter.

Fråga: Vilken kartstorlek ska man använda?

	Kartstorleken beror på hur många spelare man är och hur snart
man vill att spelet ska ta slut. Standardkartstorleken (80x50) är
tillräckligt stor för ett ganska snabbt 2-spelarspel men ger ett
*mycket* snabbt spel om > 3 spelare deltar.

	Snabba spel brukar vara otillfredställande för alla utom
vinnaren eftersom ingen har haft tid att utveckla något försvar. Om
man har > 3 spelare bör man använda en 80x80-karta. Om man är > 5
spelare bör man ha en 100x100-karta.


Fråga: Vad innebär servertillvalet "generator"?

	Den påverkar det sätt på vilket kartan skapas. Om man spelat
Freeciv några gånger utan att ändra på denna servertillvalet har
man säkerligen hört talas om (och/eller upplevt) problemen med en
alldeles för liten ö. Att behöva börja på en alldeles för liten ö kan
göra folk vansinniga. För att åtgärda detta har våra godhjärtade
hjältar till programmerare byggt in servertillvalet "generator".
- När den är satt till 1 ger det en vanlig karta med öar av olika
  (orättvisa) storlekar.
- När den är satt till 2 skapas en karta m.h.a. en pseudo-fraktal
  generator. Det innebär att berg och kullar placeras i enlighet
  med en naturlig matematisk formel.
- När den är satt till 3 skapas en lika stor ö för varje spelare,
  så att ingen kan skylla på sin ö om de förlorar.
- 0 används för färdiga kartor. Ladda en karta med /load
  /katalog/savegame.sav.gz i chatraden.

Under "generator" finns även tillvalet "startpos". Detta tillval
avgör hur många spelare som startar på samma ö. Varje "generator"-
tillval has sitt egen standardvärde som används när "startpos" är
satt till 0. Standardvärdet för "generator" 2 till exempel är 3,
vilket innbär att den försöker placera samtliga spelare på samma ö.

Fråga: Ska man förenkla spelet genom att öka mängden guld som spelarna
       får att börja med?

	Om en oerfaren spelare som spelar mot erfarna spelare föreslår
en ökning av guldmängden kommer antagligen ingen att beklaga sig.
Detta är dock inget bra sätt att lära sig att spela. Att börja med
massor av guld gör spelet mycket enklare och gör det svårare att lära
sig att hanskas med standardguldmängden. De flesta erfarna spelare
ökar inte mängden, och de vet hur de ska få mest nytta av en ökning.
Det vet inte oerfarna spelare. Därför går de i så fall samma öde till
mötes som Atlantis.

Anmärkning: Samma sak gäller inställningarna "techlevel" och
"researchspeed"

Fråga: Hur är det med de andra inställningarna?

	Resten av dem har mest att göra med vilken sorts karta som
kommer att skapas inför spelet. Att öka "specials" ger större
sannolikhet att få många tillgångar/ruta och "huts" avgör hur många
mindre stambyar det ska finnas. Att öka antalet bosättare och
utforskare gör att spelet går fortare och ökar sannolikheten att
spelare överlever barbarstammarna som i bland finns i de mindre
stambyarna.

	Inställningarna som har med järnväg att göra avgör hur mycket
en ruta ger i form av mat/sköldar/handel med järnväg och "foodbox"
bestämmer hur mycket mat varje medborgare i en stad måste ha innan en
ny person kan läggas till.

	För övrigt ger högre "mountains" mer berg, högre "deserts" ger
mer öken och så vidare.

Fråga: Hur får man en viss teknologi?

	Titta i den inbyggda hjälpen. Den visar vilka teknologier man
måste ha först.

Det går även att se detta i David Pfitzners "techtree"-karta som kan
laddas ned från <https://files.freeciv.org/contrib/charts/>.

Om det inte går man kan läsa i "data/default/techs.ruleset". Där står
vilka teknologier som man måste ha innan man kan få en given
teknologi.

Fråga: Vilka krigsenheter är bäst?

   För angrepp:

	pansar, helikopter, kryssningsmissil, slagskepp, fraktskepp,
	kärnvapen, haubits, bombflygplan.

   För försvar:

	pansar, mekaniserat infanteri, haubits, slagskepp,
	kryssningsmissil, kärnvapen.

Kom i håg att det bästa försvaret är ett kraftfullt angrepp.

Tillägg till detta dokument är välkomna!
